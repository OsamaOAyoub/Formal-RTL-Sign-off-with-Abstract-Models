package proc_states_operations;

  typedef enum { proc_states_op_Decode_2, proc_states_op_Decode_3, proc_states_op_Decode_4, proc_states_op_Decode_5, proc_states_op_Fetch_1, proc_states_op_execute_6, proc_states_op_execute_7, proc_states_op_execute_8, proc_states_op_execute_9, proc_states_op_execute_10, proc_states_op_execute_11, proc_states_op_execute_12, proc_states_op_execute_13, proc_states_op_memory_14, proc_states_op_memory_15, proc_states_op_writeback_16, proc_states_op_writeback_17, proc_states_op_writeback_18, proc_states_op_writeback_19 } proc_states_operations_t;

endpackage
