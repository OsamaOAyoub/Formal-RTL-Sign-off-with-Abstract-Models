package global_package;

  typedef bit unsigned [7:0] a_sc_unsigned_8_8[7:0];

endpackage
