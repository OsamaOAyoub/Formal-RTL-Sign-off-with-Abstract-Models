package global_package;

  const bit unsigned [31:0] CNT_SIZE = 7;

endpackage
