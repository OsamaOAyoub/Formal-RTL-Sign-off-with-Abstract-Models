package SHA512_operations;

  typedef enum { SHA512_op_DONE_9, SHA512_op_IDLE_1, SHA512_op_IDLE_2, SHA512_op_IDLE_3, SHA512_op_IDLE_4, SHA512_op_IDLE_5, SHA512_op_wait_IDLE, SHA512_op_SHARounds_8, SHA512_op_SHARounds_6, SHA512_op_SHARounds_7 } SHA512_operations_t;

endpackage
