package OptionsParser_operations;

  typedef enum { OptionsParser_op_s_DATAPARSING_14, OptionsParser_op_s_DATAPARSING_16, OptionsParser_op_s_DATAPARSING_19, OptionsParser_op_s_DATAPARSING_15, OptionsParser_op_s_DATAPARSING_17, OptionsParser_op_s_DATAPARSING_18, OptionsParser_op_s_DONE_21, OptionsParser_op_wait_s_DONE, OptionsParser_op_s_ENDPARSING_20, OptionsParser_op_s_INFOPARSING_11, OptionsParser_op_s_INFOPARSING_12, OptionsParser_op_s_INFOPARSING_9, OptionsParser_op_s_INFOPARSING_10, OptionsParser_op_s_INFOPARSING_8, OptionsParser_op_s_INFOPARSING_13, OptionsParser_op_s_READY_1, OptionsParser_op_wait_s_READY, OptionsParser_op_s_STARTPARSING_5, OptionsParser_op_s_STARTPARSING_6, OptionsParser_op_s_STARTPARSING_2, OptionsParser_op_s_STARTPARSING_3, OptionsParser_op_s_STARTPARSING_4, OptionsParser_op_s_STARTPARSING_7 } OptionsParser_operations_t;

endpackage
