package proc_states_package;

import global_package::*;


  typedef enum { IF, ID, EX, MEM, WB } e_states;

endpackage
